Accerciser
Ge ditt program en omgång hjälpmedelsfunktioner
Hjälpmedelsutforskaren Accerciser
Standardlayouten för insticksmoduler för nederpanelen
Standardlayouten för insticksmoduler för överpanelen
En lista över insticksmoduler som är inaktiverade som standard
Markeringslängd
Längden för markeringsrutan när hjälpmedelsnoder markeras
Färg för markeringsram
Färg och opacitet för markeringsramen.
Färg för markeringsfyllnad
Färg och opacitet för markeringsfyllnad.
API-bläddrare
Bläddra bland olika metoder för aktuell hjälpmedelsfunktion
Dölj privata attribut
Metod
Egenskap
Värde
IPython-konsoll
Interaktiv konsoll för manipulering av aktuell markerad hjälpmedelsfunktion
Händelseövervakare
_Övervaka händelser
Tö_m markering
Allting
Markerat program
Markerad hjälpmedelsfunktion
Källa
Händelseövervakare
Visar händelser när de inträffar från markerade typer och källor
Markera senaste händelsepost
Starta/stoppa händelseinspelning
Töm händelselogg
Antal barn
(ingen beskrivning)
Beskrivning
Tillstånd
Visa
Relationer
Attribut
_Hjälpmedelsfunktion
Genomför åtgärd
Åtgä_rd
ID
Verktygslåda
Version
_Program
Sam_ling
0, 0
Relativ position
Storlek
WIDGET
Lager
MDI-Z-ordning
Alfa
Absolut position
Ko_mponent
S_krivbord
Lokal:
_Dokument
Hyperlänk
H_ypertext
Position
Beskrivning
Lokal
_Bild
Inlo_ggningshjälpare
Markera allt
_Markering
St_römmande innehåll
Text:
Sammandrag:
Markerade kolumner
Markerade rader
Kolumner
Rader
Tabellinformation
namn (x,y)
Rubrik:
Områden:
Rad
Kolumn
Markerad cell
_Tabell
Text
Offset
Inkludera standardvärden
Start: 0
Slut: 0
Te_xt
Aktuellt värde
Minimal ökning
Maximalt värde
Minimalt värde
Vä_rde
okänd
Gränssnittsvisare
Tillåter visning av olika gränssnittsegenskaper
(inte implementerad)
Namn
URI
Start
Slut
För många valbara barn
(Redigerbar)
Snabbväljare
Insticksmodul med olika metoder för att välja hjälpmedelsfunktioner snabbt.
Inspektera senaste fokuserad hjälpmedelsfunktion
Inspektera hjälpmedelsfunktion under muspekare
Original
Dogtail
LDTP
Skripttyp
Skriptinspelare
Skapar dogtail-liknande skript
Det aktuella skriptet kommer att förloras.
Bekräfta tömning
Sche_ma:
V_alidera
Overksam
Ingen beskrivning
AT-SPI-validerare
Validerar hjälpmedel i program
Nivå
Roll
Sparar
Validerar
UNDANTAG
FEL
VARNING
INFO
FELSÖKNING
Grundläggande
Testar grundläggande hjälpmedel i grafiska program
åtgärdningsbara %s är inte fokusbar eller valbar
interaktiva %s är inte åtgärdningsbar
fler än en fokuserad widget
%s har inget textgränssnitt
%s index i förälder matchar inte barnindex
Saknar mottagare för %s-förhållande
%s saknar namn eller etikett
fokusbar %s har tabellgränssnitt, inget valgränssnittbutton has focused state without focusable state
%s har tillståndet %s utan tillståndet %s
%s tillhör inte en uppsättning
%(rolename)s index %(num)d matchar inte rad och kolumnparent indexrow and column index
%(rolename)s föräldraindex %(num1)d matchar inte rad- och kolumnindex %(num2)d
%s har inget namn eller beskrivning
_Inställningar...
_Innehåll
Accerciser kunde inte se programmen på ditt skrivbord. Du måste aktivera hjälpmedelsfunktioner för skrivbordet för att rätta till det här problemet. Vill du aktivera den nu?
Observera: Eventuella ändringar blir aktiverade efter utloggning.
